** DCIM **
** Environment setting **
.tran 0.01n 26n
.option POST
.protect
.lib "/usr/cad/cic018.l" tt
.temp 30
.unprotect
*.protect
*.lib "cic018.l" tt
*.unprotect
*********************
** Clock Parameter **
*********************
.param    CLK_Period = 2n
.param    CLK_Period_2 = 'CLK_Period/2'
.param    r_time = 1p
.param    f_time = 1p
.param    SupplyV = 1.8v
********************
* voltage setting **
********************
.global VDD GND
Vdd1 VDD 0 DC=+1.8v
Vgnd1 GND 0 DC=0v

*****************
*** My subckt ***
*****************

.subckt pFET D G S VDD
mp1 D G S VDD P_18 w=0.72u l=0.18u
.ends

.subckt nFET D G S GND
mn1 D G S GND N_18 w=0.36u l=0.18u
.ends

.subckt INV in out VDD GND
mp1	out in VDD VDD P_18 w=0.72u l=0.18u
mn1	out in GND GND N_18 w=0.36u l=0.18u
.ends

.subckt TG in C C_ out VDD GND
*Xinv1	c   c_ VDD GND INV
mp1 	out C_ in VDD P_18 w=0.72u l=0.18u
mn1	out C  in GND N_18 w=0.36u l=0.18u
.ends

.subckt DLatch_TG D C Q VDD GND
Xtg1 	D C C_ d1 VDD GND TG
Xinv1 	d1 d2 VDD GND INV
Xinv2	d2 Q  VDD GND INV
Xinv3 	C  C_ VDD GND INV
Xtg2	Q C_ C d1 VDD GND TG
.ends

.subckt W w3 w2 w1 w0 VDD GND
Xl1	GND GND w0 VDD GND DLatch_TG
Xl2	GND GND w1 VDD GND DLatch_TG
Xl3	GND GND w2 VDD GND DLatch_TG
Xl4	GND GND w3 VDD GND DLatch_TG
.ends

.subckt DLatch_tr D C Q VDD GND
Xinv1	C	C_	VDD GND INV
Xnf1	d1	C	D GND nFET
Xinv2	d1	Q_	VDD GND INV
Xinv3	Q_	Q	VDD GND INV
Xnf2	d1	C_	Q GND nFET
.ends

.subckt NOR2 in1 in2 NOR VDD GND
mp1	pd1 in1 VDD VDD P_18 w=0.72u l=0.18u
mp2	NOR in2 pd1 VDD P_18 w=0.72u l=0.18u
mn1	NOR in1 GND GND N_18 w=0.36u l=0.18u
mn2	NOR in2 GND GND N_18 w=0.36u l=0.18u
.ends

.subckt	OR2 in1 in2 OR VDD GND
Xnor	in1 in2 NOR VDD GND NOR2
Xinv	NOR OR VDD GND INV
.ends

.subckt NAND2 in1 in2 NAND VDD GND
mp1	NAND in1 VDD VDD P_18 w=0.72u l=0.18u
mp2	NAND in2 VDD VDD P_18 w=0.72u l=0.18u
mn1	NAND in1 ns1 GND N_18 w=0.36u l=0.18u
mn2	ns1  in2 GND GND N_18 w=0.36u l=0.18u
.ends

.subckt AND2 in1 in2 AND VDD GND
Xnand	in1 in2 NAND VDD GND NAND2
Xinv	NAND	AND VDD GND INV
.ends

*** XNOR ***
.subckt XNOR2 A B XNOR VDD GND
Xinv1	A A_ VDD GND INV
Xinv2	B B_ VDD GND INV
Xnand1	A  B ndAB VDD GND NAND2
Xor1	A  B AorB VDD GND OR2
Xnand2	ndAB AorB XNOR VDD GND NAND2
.ends
*** XOR ***
.subckt XOR2 A B XOR VDD GND
Xxnor	A B XNOR VDD GND XNOR2
Xinv1	XNOR XOR VDD GND INV
.ends
*** Half Adder ***
.subckt HalfAdd1 A B Cout Sum VDD GND
Xxor	A B Sum  VDD GND XOR2
Xand	A B Cout VDD GND AND2
.ends
*** Full Adder ***
.subckt FullAdd1 A B C Cout S VDD GND
mp1  x1  A VDD VDD P_18 w=0.72u l=0.18u
mp2  x1  B VDD VDD P_18 w=0.72u l=0.18u
mp3  x3  A VDD VDD P_18 w=0.72u l=0.18u
mp4  cob B x3  VDD P_18 w=0.72u l=0.18u
mp5  cob C x1  VDD P_18 w=0.72u l=0.18u

mn1  cob C x2  GND N_18 w=0.36u l=0.18u
mn2  x2  A GND GND N_18 w=0.36u l=0.18u
mn3  x2  B GND GND N_18 w=0.36u l=0.18u
mn4  cob B x4  GND N_18 w=0.36u l=0.18u 
mn5  x4  A GND GND N_18 w=0.36u l=0.18u 

mp6 x5  A VDD VDD P_18 w=0.72u l=0.18u 
mp7 x5  B VDD VDD P_18 w=0.72u l=0.18u 
mp8 x5  C VDD VDD P_18 w=0.72u l=0.18u 
mp9 sb  cob x5 VDD P_18 w=0.72u l=0.18u 

mn6 sb cob x6 GND N_18 w=0.36u l=0.18u 
mn7 x6 A GND GND N_18 w=0.36u l=0.18u 
mn8 x6 B GND GND N_18 w=0.36u l=0.18u 
mn9 x6 C GND GND N_18 w=0.36u l=0.18u

mp10 Cout cob VDD VDD P_18 w=0.72u l=0.18u
mn10 Cout cob GND GND N_18 w=0.36u l=0.18u

mp11 x7 A VDD VDD P_18 w=0.72u l=0.18u 
mp12 x8 B x7  VDD P_18 w=0.72u l=0.18u 
mp13 sb C x8  VDD P_18 w=0.72u l=0.18u

mn11 sb C  x9  GND N_18 w=0.36u l=0.18u 
mn12 x9 B  x10 GND N_18 w=0.36u l=0.18u 
mn13 x10 A GND GND N_18 w=0.36u l=0.18u 

mp14 S sb VDD VDD P_18 w=0.72u l=0.18u 
mn14 S sb GND GND N_18 w=0.36u l=0.18u 
.ends

*** Full Adder 4 bits ***
.subckt FullAdd4 A3 A2 A1 A0 B3 B2 B1 B0 Cin S4 S3 S2 S1 S0 VDD GND
Xfa1	A0 B0 Cin C0 S0 VDD GND FullAdd1
Xfa2	A1 B1 C0  C1 S1 VDD GND FullAdd1
Xfa3	A2 B2 C1  C2 S2 VDD GND FullAdd1
Xfa4	A3 B3 C2  S4 S3 VDD GND FullAdd1
.ends
*** Full Adder 5 bits ***
.subckt FullAdd5 A4 A3 A2 A1 A0 B4 B3 B2 B1 B0 Cin S5 S4 S3 S2 S1 S0 VDD GND
Xfa4b	A3 A2 A1 A0 B3 B2 B1 B0 Cin C3 S3 S2 S1 S0 VDD GND FullAdd4
Xfa5	A4 B4 C3 S5 S4 VDD GND FullAdd1
.ends
*** Full Adder 10 bits ***
.subckt FullAdd10 A9 A8 A7 A6 A5 A4 A3 A2 A1 A0 B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 Cin S10 S9 S8 S7 S6 S5 S4 S3 S2 S1 S0 VDD GND
Xfa5b1	A4 A3 A2 A1 A0 B4 B3 B2 B1 B0 Cin C4 S4 S3 S2 S1 S0 VDD GND FullAdd5
Xfa5b2	A9 A8 A7 A6 A5 B9 B8 B7 B6 B5 C4 S10 S9 S8 S7 S6 S5 VDD GND FullAdd5
.ends

.subckt FullAdd10b A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 B0 B1 B2 B3 B4 B5 B6 B7 B8 B9 Cin S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 VDD GND
Xfa5b1	A4 A3 A2 A1 A0 B4 B3 B2 B1 B0 Cin C4 S4 S3 S2 S1 S0 VDD GND FullAdd5
Xfa5b2	A9 A8 A7 A6 A5 B9 B8 B7 B6 B5 C4 S10 S9 S8 S7 S6 S5 VDD GND FullAdd5
.ends

*** Flip Flop ***
.subckt DFF D CLK Q VDD GND
Xinv 	CLK CLK_ VDD GND INV
Xdl1	D CLK_ Y VDD GND DLatch_TG
Xdl2	Y CLK  Q VDD GND DLatch_TG
.ends

******************
*** End subckt ***
******************
**********************************************
*** Don't modify the pin name in this file ***
**********************************************
Xdcim I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O10 O11 O12 O13 O14 O15 O16 O17 O18 O19 O20 O21 O22 O23 O24 O25 O26 O27 O28 O29 O30 O31 O32 O33 O34 O35 O36 O37 O38 O39 O40 O41 O42 O43 O44 O45 O46 O47 O48 O49 O50 O51 O52 O53 O54 O55 O56 O57 O58 O59 O60 O61 O62 O63 O64 O65 O66 O67 O68 O69 O70 O71 O72 O73 O74 O75 O76 O77 O78 O79 O80 O81 O82 O83 O84 O85 O86 O87 O88 O89 O90 O91 O92 O93 O94 O95 O96 O97 O98 O99 O100 O101 O102 O103 O104 O105 O106 O107 O108 O109 O110 O111 O112 O113 O114 O115 O116 O117 O118 O119 O120 O121 O122 O123 O124 O125 O126 O127 O128 O129 O130 O131 O132 O133 O134 O135 O136 O137 O138 O139 O140 O141 O142 O143 O144 O145 O146 O147 O148 O149 O150 O151 O152 O153 O154 O155 O156 O157 O158 O159 O160 O161 O162 O163 O164 O165 O166 O167 O168 O169 OUT_VAL DCIM

*** Initial Condition ***
*** Initial Weights column 1
.ic V(Xdcim.Xw1.w3)=0v V(Xdcim.Xw1.w2)=0v V(Xdcim.Xw1.w1)=0v V(Xdcim.Xw1.w0)=0v
.ic V(Xdcim.Xw2.w3)=0v V(Xdcim.Xw2.w2)=0v V(Xdcim.Xw2.w1)=0v V(Xdcim.Xw2.w0)=1.8v
.ic V(Xdcim.Xw3.w3)=0v V(Xdcim.Xw3.w2)=0v V(Xdcim.Xw3.w1)=1.8v V(Xdcim.Xw3.w0)=0v
.ic V(Xdcim.Xw4.w3)=0v V(Xdcim.Xw4.w2)=0v V(Xdcim.Xw4.w1)=1.8v V(Xdcim.Xw4.w0)=1.8v
.ic V(Xdcim.Xw5.w3)=0v V(Xdcim.Xw5.w2)=1.8v V(Xdcim.Xw5.w1)=0v V(Xdcim.Xw5.w0)=0v
.ic V(Xdcim.Xw6.w3)=0v V(Xdcim.Xw6.w2)=1.8v V(Xdcim.Xw6.w1)=0v V(Xdcim.Xw6.w0)=1.8v
.ic V(Xdcim.Xw7.w3)=0v V(Xdcim.Xw7.w2)=1.8v V(Xdcim.Xw7.w1)=1.8v V(Xdcim.Xw7.w0)=0v
.ic V(Xdcim.Xw8.w3)=0v V(Xdcim.Xw8.w2)=1.8v V(Xdcim.Xw8.w1)=1.8v V(Xdcim.Xw8.w0)=1.8v
.ic V(Xdcim.Xw9.w3)=1.8v V(Xdcim.Xw9.w2)=0v V(Xdcim.Xw9.w1)=0v V(Xdcim.Xw9.w0)=0v
.ic V(Xdcim.Xw10.w3)=1.8v V(Xdcim.Xw10.w2)=0v V(Xdcim.Xw10.w1)=0v V(Xdcim.Xw10.w0)=1.8v
.ic V(Xdcim.Xw11.w3)=1.8v V(Xdcim.Xw11.w2)=0v V(Xdcim.Xw11.w1)=1.8v V(Xdcim.Xw11.w0)=0v
.ic V(Xdcim.Xw12.w3)=1.8v V(Xdcim.Xw12.w2)=0v V(Xdcim.Xw12.w1)=1.8v V(Xdcim.Xw12.w0)=1.8v
.ic V(Xdcim.Xw13.w3)=1.8v V(Xdcim.Xw13.w2)=1.8v V(Xdcim.Xw13.w1)=0v V(Xdcim.Xw13.w0)=0v
.ic V(Xdcim.Xw14.w3)=1.8v V(Xdcim.Xw14.w2)=1.8v V(Xdcim.Xw14.w1)=0v V(Xdcim.Xw14.w0)=1.8v
.ic V(Xdcim.Xw15.w3)=1.8v V(Xdcim.Xw15.w2)=1.8v V(Xdcim.Xw15.w1)=1.8v V(Xdcim.Xw15.w0)=0v
.ic V(Xdcim.Xw16.w3)=1.8v V(Xdcim.Xw16.w2)=1.8v V(Xdcim.Xw16.w1)=1.8v V(Xdcim.Xw16.w0)=1.8v

*************************

.subckt DCIM I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O10 O11 O12 O13 O14 O15 O16 O17 O18 O19 O20 O21 O22 O23 O24 O25 O26 O27 O28 O29 O30 O31 O32 O33 O34 O35 O36 O37 O38 O39 O40 O41 O42 O43 O44 O45 O46 O47 O48 O49 O50 O51 O52 O53 O54 O55 O56 O57 O58 O59 O60 O61 O62 O63 O64 O65 O66 O67 O68 O69 O70 O71 O72 O73 O74 O75 O76 O77 O78 O79 O80 O81 O82 O83 O84 O85 O86 O87 O88 O89 O90 O91 O92 O93 O94 O95 O96 O97 O98 O99 O100 O101 O102 O103 O104 O105 O106 O107 O108 O109 O110 O111 O112 O113 O114 O115 O116 O117 O118 O119 O120 O121 O122 O123 O124 O125 O126 O127 O128 O129 O130 O131 O132 O133 O134 O135 O136 O137 O138 O139 O140 O141 O142 O143 O144 O145 O146 O147 O148 O149 O150 O151 O152 O153 O154 O155 O156 O157 O158 O159 O160 O161 O162 O163 O164 O165 O166 O167 O168 O169 OUT_VAL

*** Weight ***
Xw1	W13 W12 W11 W10 VDD GND W
Xw2	W23 W22 W21 W20 VDD GND W
Xw3	W33 W32 W31 W30 VDD GND W
Xw4	W43 W42 W41 W40 VDD GND W
Xw5	W53 W52 W51 W50 VDD GND W
Xw6	W63 W62 W61 W60 VDD GND W
Xw7	W73 W72 W71 W70 VDD GND W
Xw8	W83 W82 W81 W80 VDD GND W
Xw9	W93 W92 W91 W90 VDD GND W
Xw10	W103 W102 W101 W100 VDD GND W
Xw11	W113 W112 W111 W110 VDD GND W
Xw12	W123 W122 W121 W120 VDD GND W
Xw13	W133 W132 W131 W130 VDD GND W
Xw14	W143 W142 W141 W140 VDD GND W
Xw15	W153 W152 W151 W150 VDD GND W
Xw16	W163 W162 W161 W160 VDD GND W
**************

Xdcim11 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O10 O11 O12 O13 O14 O15 O16 O17 O18 O19 O20 O21 O22 O23 O24 O25 O26 O27 O28 O29 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM32_2

Xdcim22 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O30 O31 O32 O33 O34 O35 O36 O37 O38 O39 O40 O41 O42 O43 O44 O45 O46 O47 O48 O49 OUT_VAL W33 W32 W31 W30 W43 W42 W41 W40 DCIM32_2

Xdcim33 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O50 O51 O52 O53 O54 O55 O56 O57 O58 O59 O60 O61 O62 O63 O64 O65 O66 O67 O68 O69 OUT_VAL W53 W52 W51 W50 W63 W62 W61 W60 DCIM32_2

Xdcim44 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O70 O71 O72 O73 O74 O75 O76 O77 O78 O79 O80 O81 O82 O83 O84 O85 O86 O87 O88 O89 OUT_VAL W73 W72 W71 W70 W83 W82 W81 W80 DCIM32_2

Xdcim55 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O90 O91 O92 O93 O94 O95 O96 O97 O98 O99 O100 O101 O102 O103 O104 O105 O106 O107 O108 O109 OUT_VAL W93 W92 W91 W90 W103 W102 W101 W100 DCIM32_2

Xdcim66 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O110 O111 O112 O113 O114 O115 O116 O117 O118 O119 O120 O121 O122 O123 O124 O125 O126 O127 O128 O129 OUT_VAL W113 W112 W111 W110 W123 W122 W121 W120 DCIM32_2

Xdcim77 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O130 O131 O132 O133 O134 O135 O136 O137 O138 O139 O140 O141 O142 O143 O144 O145 O146 O147 O148 O149 OUT_VAL W133 W132 W131 W130 W143 W142 W141 W140 DCIM32_2

Xdcim88 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O150 O151 O152 O153 O154 O155 O156 O157 O158 O159 O160 O161 O162 O163 O164 O165 O166 O167 O168 O169 OUT_VAL W153 W152 W151 W150 W163 W162 W161 W160 DCIM32_2

.ends
*****************
*** call cell ***
*****************
.subckt DCIM32_2 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31 I32 IN_VAL CLK RST O10 O11 O12 O13 O14 O15 O16 O17 O18 O19 O20 O21 O22 O23 O24 O25 O26 O27 O28 O29 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20
Xdcim1 I1 I2 I3 I4 IN_VAL CLK RST p110 p111 p112 p113 p114 p115 p116 p117 p118 p119 p120 p121 p122 p123 p124 p125 p126 p127 p128 p129 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2
Xdcim2 I5 I6 I7 I8 IN_VAL CLK RST p210 p211 p212 p213 p214 p215 p216 p217 p218 p219 p220 p221 p222 p223 p224 p225 p226 p227 p228 p229 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2

Xdcim3 I9 I10 I11 I12 IN_VAL CLK RST p310 p311 p312 p313 p314 p315 p316 p317 p318 p319 p320 p321 p322 p323 p324 p325 p326 p327 p328 p329 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2
Xdcim4 I13 I14 I15 I16 IN_VAL CLK RST p410 p411 p412 p413 p414 p415 p416 p417 p418 p419 p420 p421 p422 p423 p424 p425 p426 p427 p428 p429 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2

Xdcim5 I17 I18 I19 I20 IN_VAL CLK RST p510 p511 p512 p513 p514 p515 p516 p517 p518 p519 p520 p521 p522 p523 p524 p525 p526 p527 p528 p529 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2
Xdcim6 I21 I22 I23 I24 IN_VAL CLK RST p610 p611 p612 p613 p614 p615 p616 p617 p618 p619 p620 p621 p622 p623 p624 p625 p626 p627 p628 p629 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2

Xdcim7 I25 I26 I27 I28 IN_VAL CLK RST p710 p711 p712 p713 p714 p715 p716 p717 p718 p719 p720 p721 p722 p723 p724 p725 p726 p727 p728 p729 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2
Xdcim8 I29 I30 I31 I32 IN_VAL CLK RST p810 p811 p812 p813 p814 p815 p816 p817 p818 p819 p820 p821 p822 p823 p824 p825 p826 p827 p828 p829 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20 DCIM4_2
*** Col 1
Xfa1	p110 p111 p112 p113 p114 p115 p116 p117 p118 p119 p210 p211 p212 p213 p214 p215 p216 p217 p218 p219 GND a0 a1 a2 a3 a4 a5 a6 a7 a8 a9 a10 VDD GND FullAdd10b
Xfa2 	p310 p311 p312 p313 p314 p315 p316 p317 p318 p319 p410 p411 p412 p413 p414 p415 p416 p417 p418 p419 GND b0 b1 b2 b3 b4 b5 b6 b7 b8 b9 b10 VDD GND FullAdd10b
Xfa3	p510 p511 p512 p513 p514 p515 p516 p517 p518 p519 p610 p611 p612 p613 p614 p615 p616 p617 p618 p619 GND c0 c1 c2 c3 c4 c5 c6 c7 c8 c9 c10 VDD GND FullAdd10b
Xfa4	p710 p711 p712 p713 p714 p715 p716 p717 p718 p719 p810 p811 p812 p813 p814 p815 p816 p817 p818 p819 GND d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 d10 VDD GND FullAdd10b

Xfa5	a0 a1 a2 a3 a4 a5 a6 a7 a8 a9 b0 b1 b2 b3 b4 b5 b6 b7 b8 b9 GND e0 e1 e2 e3 e4 e5 e6 e7 e8 e9 e10 VDD GND FullAdd10b
Xfa6	c0 c1 c2 c3 c4 c5 c6 c7 c8 c9 d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 GND f0 f1 f2 f3 f4 f5 f6 f7 f8 f9 f10 VDD GND FullAdd10b

Xfa7	e0 e1 e2 e3 e4 e5 e6 e7 e8 e9 f0 f1 f2 f3 f4 f5 f6 f7 f8 f9 GND O10 O11 O12 O13 O14 O15 O16 O17 O18 O19 Ox VDD GND FullAdd10b
*** Col 2
Xfa8	p120 p121 p122 p123 p124 p125 p126 p127 p128 p129 p220 p221 p222 p223 p224 p225 p226 p227 p228 p229 GND g0 g1 g2 g3 g4 g5 g6 g7 g8 g9 g10 VDD GND FullAdd10b
Xfa9 	p320 p321 p322 p323 p324 p325 p326 p327 p328 p329 p420 p421 p422 p423 p424 p425 p426 p427 p428 p429 GND h0 h1 h2 h3 h4 h5 h6 h7 h8 h9 h10 VDD GND FullAdd10b
Xfa10	p520 p521 p522 p523 p524 p525 p526 p527 p528 p529 p620 p621 p622 p623 p624 p625 p626 p627 p628 p629 GND i0 i1 i2 i3 i4 i5 i6 i7 i8 i9 i10 VDD GND FullAdd10b
Xfa11	p720 p721 p722 p723 p724 p725 p726 p727 p728 p729 p820 p821 p822 p823 p824 p825 p826 p827 p828 p829 GND j0 j1 j2 j3 j4 j5 j6 j7 j8 j9 j10 VDD GND FullAdd10b

Xfa12	g0 g1 g2 g3 g4 g5 g6 g7 g8 g9 h0 h1 h2 h3 h4 h5 h6 h7 h8 h9 GND k0 k1 k2 k3 k4 k5 k6 k7 k8 k9 k10 VDD GND FullAdd10b
Xfa13	i0 i1 i2 i3 i4 i5 i6 i7 i8 i9 j0 j1 j2 j3 j4 j5 j6 j7 j8 j9 GND l0 l1 l2 l3 l4 l5 l6 l7 l8 l9 l10 VDD GND FullAdd10b

Xfa14	k0 k1 k2 k3 k4 k5 k6 k7 k8 k9 l0 l1 l2 l3 l4 l5 l6 l7 l8 l9 GND O20 O21 O22 O23 O24 O25 O26 O27 O28 O29 Ox VDD GND FullAdd10b
.ends

******************
*** DCIM block ***
******************
.subckt DCIM4_2 I1 I2 I3 I4 IN_VAL CLK RST O10 O11 O12 O13 O14 O15 O16 O17 O18 O19 O20 O21 O22 O23 O24 O25 O26 O27 O28 O29 OUT_VAL W13 W12 W11 W10 W23 W22 W21 W20
*** Inverse CLK
Xinv0 CLK CLK_ VDD GND INV
*** Input rounds
** Col 1
Xiw11	ii1 W13 W12 W11 W10 o113 o112 o111 o110 VDD GND IdotW
Xiw12	ii2 W13 W12 W11 W10 o123 o122 o121 o120 VDD GND IdotW
Xiw13	ii3 W13 W12 W11 W10 o133 o132 o131 o130 VDD GND IdotW
Xiw14	ii4 W13 W12 W11 W10 o143 o142 o141 o140 VDD GND IdotW
** Col 2
Xiw21	ii1 W23 W22 W21 W20 o213 o212 o211 o210 VDD GND IdotW
Xiw22	ii2 W23 W22 W21 W20 o223 o222 o221 o220 VDD GND IdotW
Xiw23	ii3 W23 W22 W21 W20 o233 o232 o231 o230 VDD GND IdotW
Xiw24	ii4 W23 W22 W21 W20 o243 o242 o241 o240 VDD GND IdotW
*** Adder Tree ***
** Add Col 1 
* I1 I2
Xfa4b1	o113 o112 o111 o110 o123 o122 o121 o120 GND i12_4 i12_3 i12_2 i12_1 i12_0 VDD GND FullAdd4
* I3 I4
Xfa4b2	o133 o132 o131 o130 o143 o142 o141 o140 GND i34_4 i34_3 i34_2 i34_1 i34_0 VDD GND FullAdd4
* 5 bits part
Xfa5b1	i12_4 i12_3 i12_2 i12_1 i12_0 i34_4 i34_3 i34_2 i34_1 i34_0 GND c1_5 c1_4 c1_3 c1_2 c1_1 c1_0 VDD GND FullAdd5

* To 10 bits full adder and cycle with register and shift
Xfa9b1	GND GND GND GND c1_5 c1_4 c1_3 c1_2 c1_1 c1_0 O18 O17 O16 O15 O14 O13 O12 O11 O10 GND GND Px P19 P18 P17 P16 P15 P14 P13 P12 P11 P10 VDD GND FullAdd10
* add into register
*Xrg10	fa19 fa18 fa17 fa16 fa15 fa14 fa13 fa12 fa11 fa10 CLK VDD P19 P18 P17 P16 P15 P14 P13 P12 P11 P10 VDD GND Register10
* Register to Shift
*Xrg11	P18 P17 P16 P15 P14 P13 P12 P11 P10 GND CLK_ RST sh19 sh18 sh17 sh16 sh15 sh14 sh13 sh12 sh11 sh10 VDD GND Register10

** Add Col 2
* I1 I2 
Xfa4b3	o213 o212 o211 o210 o223 o222 o221 o220 GND i212_4 i212_3 i212_2 i212_1 i212_0 VDD GND FullAdd4
* I3 I4
Xfa4b4 	o233 o232 o231 o230 o243 o242 o241 o240 GND i234_4 i234_3 i234_2 i234_1 i234_0 VDD GND FullAdd4
* 5 bits part
Xfa5b2	i212_4 i212_3 i212_2 i212_1 i212_0 i234_4 i234_3 i234_2 i234_1 i234_0 GND c2_5 c2_4 c2_3 c2_2 c2_1 c2_0 VDD GND FullAdd5
* Add and put into output register
Xfa9b2  GND GND GND GND c2_5 c2_4 c2_3 c2_2 c2_1 c2_0 O28 O27 O26 O25 O24 O23 O22 O21 O20 GND GND Py P29 P28 P27 P26 P25 P24 P23 P22 P21 P20 VDD GND FullAdd10

*** OUT_VAL == 1
Xoutnow IN_VAL CLK OUT_VAL VDD GND OUT_NOW

Xcontrol_in I1 I2 I3 I4 CLK IN_VAL ii1 ii2 ii3 ii4 CON_IN
Xcontrol_out1 P10 P11 P12 P13 P14 P15 P16 P17 P18 P19 CLK RST O10 O11 O12 O13 O14 O15 O16 O17 O18 O19 CON_OUT
Xcontrol_out2 P20 P21 P22 P23 P24 P25 P26 P27 P28 P29 CLK RST O20 O21 O22 O23 O24 O25 O26 O27 O28 O29 CON_OUT
.ends

************************
*** input controller ***
************************
.subckt CON_IN I1 I2 I3 I4 CLK IN_VAL ii1 ii2 ii3 ii4
Xand1 I1 IN_VAL out1 VDD GND AND2
Xand2 I2 IN_VAL out2 VDD GND AND2
Xand3 I3 IN_VAL out3 VDD GND AND2
Xand4 I4 IN_VAL out4 VDD GND AND2
Xff1  out1 CLK ii1 VDD GND DFF
Xff2  out2 CLK ii2 VDD GND DFF
Xff3  out3 CLK ii3 VDD GND DFF
Xff4  out4 CLK ii4 VDD GND DFF
*** Your code ***
.ends
*** Add round subcircuit
.subckt IdotW ii w3 w2 w1 w0 o3 o2 o1 o0 VDD GND
Xand1 ii w0 o0 VDD GND AND2
Xand2 ii w1 o1 VDD GND AND2
Xand3 ii w2 o2 VDD GND AND2
Xand4 ii w3 o3 VDD GND AND2
.ends
*************************
*** output controller ***
*************************
.subckt OUT_NOW IN_VAL CLK OUT_VAL VDD GND
Xff1	IN_VAL CLK    Pre_in   VDD GND DFF
Xinv	IN_VAL IN_bar	       VDD GND INV
Xand	Pre_in IN_bar Fall     VDD GND AND2
Xff2	Fall   CLK    OUT_VAL  VDD GND DFF
.ends

.subckt CON_OUT P0 P1 P2 P3 P4 P5 P6 P7 P8 P9 CLK RST O0 O1 O2 O3 O4 O5 O6 O7 O8 O9 
Xand0	P0 RST P00 VDD GND AND2
Xand1   P1 RST P11 VDD GND AND2
Xand2   P2 RST P22 VDD GND AND2
Xand3   P3 RST P33 VDD GND AND2
Xand4   P4 RST P44 VDD GND AND2
Xand5   P5 RST P55 VDD GND AND2
Xand6   P6 RST P66 VDD GND AND2
Xand7   P7 RST P77 VDD GND AND2
Xand8   P8 RST P88 VDD GND AND2
Xand9   P9 RST P99 VDD GND AND2
Xff0	P00 CLK O0 VDD GND DFF
Xff1    P11 CLK O1 VDD GND DFF
Xff2    P22 CLK O2 VDD GND DFF
Xff3    P33 CLK O3 VDD GND DFF
Xff4    P44 CLK O4 VDD GND DFF
Xff5    P55 CLK O5 VDD GND DFF
Xff6    P66 CLK O6 VDD GND DFF
Xff7    P77 CLK O7 VDD GND DFF
Xff8    P88 CLK O8 VDD GND DFF
Xff9    P99 CLK O9 VDD GND DFF
.ends

**************************
*** Simulation setting ***
**************************
Vclk CLK 0 PULSE(0v SupplyV 0 r_time f_time CLK_Period_2 CLK_Period)

Vrst RST 0 PWL 0n SupplyV
+ 'CLK_Period*1.5' SupplyV 'CLK_Period*1.5+f_time' 0v 'CLK_Period*2.5' 0v 'CLK_Period*2.5+r_time' SupplyV
+ 'CLK_Period*6.5' SupplyV 'CLK_Period*6.5+f_time' 0v 'CLK_Period*7.5' 0v 'CLK_Period*7.5+r_time' SupplyV

Vval IN_VAL 0 PWL 0n 0v
+ 'CLK_Period*1' 0v 'CLK_Period*1+f_time' SupplyV 'CLK_Period*5' SupplyV 'CLK_Period*5+r_time' 0v
+ 'CLK_Period*6' 0v 'CLK_Period*6+f_time' SupplyV 'CLK_Period*10' SupplyV 'CLK_Period*10+r_time' 0v

*8 -> 15
VD1 I1 0 PWL 0n 0v
+ 'CLK_Period*1' 0v 'CLK_Period*1+r_time' SupplyV 'CLK_Period*2' SupplyV 'CLK_Period*2+f_time' 0v
+ 'CLK_Period*6' 0v 'CLK_Period*6+r_time' SupplyV 'CLK_Period*10' SupplyV 'CLK_Period*10+f_time' 0v
*2 -> 14
VD2 I2 0 PWL 0n 0v
+ 'CLK_Period*3' 0v 'CLK_Period*3+r_time' SupplyV 'CLK_Period*4' SupplyV 'CLK_Period*4+r_time' 0v
+ 'CLK_Period*6' 0v 'CLK_Period*6+r_time' SupplyV 'CLK_Period*9' SupplyV 'CLK_Period*9+f_time' 0v
*3 -> 13
VD3 I3 0 PWL 0n 0v
+ 'CLK_Period*3' 0v 'CLK_Period*3+r_time' SupplyV 'CLK_Period*5' SupplyV 'CLK_Period*5+f_time' 0v
+ 'CLK_Period*6' 0v 'CLK_Period*6+r_time' SupplyV 'CLK_Period*8' SupplyV 'CLK_Period*8+f_time' 0v
+ 'CLK_Period*9' 0v 'CLK_Period*9+r_time' SupplyV 'CLK_Period*10' SupplyV 'CLK_Period*10+f_time' 0v
*7 -> 12
VD4 I4 0 PWL 0n 0v
+ 'CLK_Period*2' 0v 'CLK_Period*2+r_time' SupplyV 'CLK_Period*5' SupplyV 'CLK_Period*5+r_time' 0v
+ 'CLK_Period*6' 0v 'CLK_Period*6+r_time' SupplyV 'CLK_Period*8' SupplyV 'CLK_Period*8+f_time' 0v

*******************
*** Measurement ***
*******************
.measure TRAN td
+ TRIG V(Xdcim.ii1) VAL=0.9 RISE=1
+ TARG V(Xdcim.P10)  VAL=0.9 RISE=1

.measure TRAN pwr AVG POWER
