* File: /home/VLSI_1131/tsx1136010/hw02/spice/post_sim/hw2/XOR3_pex/XOR3_pex.cir
* Created: Sat Nov 16 21:15:46 2024
* Program "Calibre xRC"
* Version "v2020.2_14.12"
* 
.include "/home/VLSI_1131/tsx1136010/hw02/spice/post_sim/hw2/XOR3_pex/XOR3_pex.cir.pex"
.subckt XOR3  A B GND VDD C S
* 
* S	S
* C	C
* VDD	VDD
* GND	GND
* B	B
* A	A
M0 N_2_M0_d N_A_M0_g N_GND_M0_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07 AD=2.968e-13
+ AS=2.968e-13 PD=1.65e-06 PS=1.65e-06
M1 N_GND_M1_d N_A_M1_g N_3_M1_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07
+ AD=1.5105e-13 AS=3.127e-13 PD=5.7e-07 PS=1.71e-06
M2 N_6_M2_d N_2_M2_g N_GND_M2_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07 AD=3.074e-13
+ AS=1.5105e-13 PD=1.69e-06 PS=5.7e-07
M3 N_14_M3_d N_B_M3_g N_GND_M3_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07
+ AD=2.915e-13 AS=3.021e-13 PD=1.63e-06 PS=1.67e-06
M4 N_3_M4_d N_14_M4_g N_10_M4_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07
+ AD=1.5105e-13 AS=3.127e-13 PD=5.7e-07 PS=1.71e-06
M5 N_13_M5_d N_B_M5_g N_3_M5_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07 AD=3.074e-13
+ AS=1.5105e-13 PD=1.69e-06 PS=5.7e-07
M6 N_6_M6_d N_B_M6_g N_10_M6_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07 AD=1.5105e-13
+ AS=3.127e-13 PD=5.7e-07 PS=1.71e-06
M7 N_13_M7_d N_14_M7_g N_6_M7_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07 AD=3.074e-13
+ AS=1.5105e-13 PD=1.69e-06 PS=5.7e-07
M8 N_16_M8_d N_C_M8_g N_GND_M8_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07
+ AD=2.968e-13 AS=2.968e-13 PD=1.65e-06 PS=1.65e-06
M9 N_S_M9_d N_16_M9_g N_13_M9_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07
+ AD=1.5105e-13 AS=3.127e-13 PD=5.7e-07 PS=1.71e-06
M10 N_10_M10_d N_C_M10_g N_S_M10_s N_GND_M0_b N_18 L=1.8e-07 W=5.3e-07
+ AD=3.074e-13 AS=1.5105e-13 PD=1.69e-06 PS=5.7e-07
M11 N_2_M11_d N_A_M11_g N_VDD_M11_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=6.72e-13 AS=6.72e-13 PD=2.32e-06 PS=2.32e-06
M12 N_VDD_M12_d N_A_M12_g N_4_M12_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.42e-13 AS=6.96e-13 PD=5.7e-07 PS=2.36e-06
M13 N_5_M13_d N_2_M13_g N_VDD_M13_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=7.2e-13 AS=3.42e-13 PD=2.4e-06 PS=5.7e-07
M14 N_14_M14_d N_B_M14_g N_VDD_M14_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=6.72e-13 AS=6.72e-13 PD=2.32e-06 PS=2.32e-06
M15 N_4_M15_d N_14_M15_g N_11_M15_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.42e-13 AS=6.96e-13 PD=5.7e-07 PS=2.36e-06
M16 N_12_M16_d N_B_M16_g N_4_M16_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=7.2e-13 AS=3.42e-13 PD=2.4e-06 PS=5.7e-07
M17 N_5_M17_d N_B_M17_g N_11_M17_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.42e-13 AS=6.96e-13 PD=5.7e-07 PS=2.36e-06
M18 N_12_M18_d N_14_M18_g N_5_M18_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=7.2e-13 AS=3.42e-13 PD=2.4e-06 PS=5.7e-07
M19 N_16_M19_d N_C_M19_g N_VDD_M19_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=6.72e-13 AS=6.72e-13 PD=2.32e-06 PS=2.32e-06
M20 N_S_M20_d N_16_M20_g N_12_M20_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.42e-13 AS=6.96e-13 PD=5.7e-07 PS=2.36e-06
M21 N_11_M21_d N_C_M21_g N_S_M21_s N_VDD_M11_b P_18 L=1.8e-07 W=1.2e-06
+ AD=7.2e-13 AS=3.42e-13 PD=2.4e-06 PS=5.7e-07
*
.include "/home/VLSI_1131/tsx1136010/hw02/spice/post_sim/hw2/XOR3_pex/XOR3_pex.cir.XOR3.pxi"
*
.ends
*
*
